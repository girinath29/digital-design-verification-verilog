module not_gate_df (
    input  wire a,
    output wire y
);
    assign y = ~a;
endmodule
