module or_gate_str (
    input  wire a,
    input  wire b,
    output wire y
);
    or u1 (y, a, b);
endmodule
