module not_gate_str (
    input  wire a,
    output wire y
);
    not u1 (y, a);
endmodule
