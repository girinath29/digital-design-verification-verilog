module and_gate_str (
    input  wire a,
    input  wire b,
    output wire y
);
    and u1 (y, a, b);
endmodule
