module nand_gate_df (
    input  wire a,
    input  wire b,
    output wire y
);
    assign y = ~(a & b);
endmodule
